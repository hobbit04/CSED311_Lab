module calculate_next_state(
    input [3:0] added_state,  // state + 1
    input [6:0] opcode,
    input [3:0] AddrCtrl,
    output reg [3:0] next_state
);
    
    always @(*) begin
        
    end
endmodule